LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

ENTITY DADO IS PORT(
    CLK, CLR, PARO : IN STD_LOGIC;
    DISPLAY:INOUT STD_LOGIC_VECTOR(6 DOWNTO 0)

);
END ENTITY DADO;

ARCHITECTURE A_DADO OF DADO IS
TYPE ESTADOS IS (A,B,C,D,E,F,APAGADO);
SIGNAL EDO_PRE, EDO_FUT: ESTADOS;
CONSTANT DIG1:STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001111";
CONSTANT DIG2:STD_LOGIC_VECTOR(6 DOWNTO 0):= "0010010";
CONSTANT DIG3:STD_LOGIC_VECTOR(6 DOWNTO 0):= "0000110";
CONSTANT DIG4:STD_LOGIC_VECTOR(6 DOWNTO 0):= "1001100";
CONSTANT DIG5:STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100100";
CONSTANT DIG6:STD_LOGIC_VECTOR(6 DOWNTO 0):= "0100000";
SIGNAL CONTADOR: UNSIGNED(31 DOWNTO 0):= (OTHERS=>'0');
SIGNAL DIV_CLK: STD_LOGIC:='0';
CONSTANT DIVISOR: INTEGER:= 2700000;


BEGIN 
PROCESS(CLK)IS
BEGIN
    IF RISING_EDGE(CLK)THEN
        IF CONTADOR>=TO_UNSIGNED(DIVISOR,32)THEN
            CONTADOR<=(OTHERS=>'0');
            DIV_CLK<=NOT DIV_CLK;
        ELSE
            CONTADOR<= CONTADOR + 1;
        END IF;
    END IF;
END PROCESS;

DIAGRAMA:PROCESS(EDO_PRE, PARO) IS
BEGIN
CASE EDO_PRE IS

    WHEN A=>DISPLAY<=DIG1;
        IF (PARO='0') THEN
            EDO_FUT<=B;
        ELSE
            EDO_FUT<=A;
        END IF;

WHEN B=>DISPLAY<=DIG2;
        IF (PARO='0') THEN
            EDO_FUT<=C;
        ELSE
            EDO_FUT<=B;
        END IF;

WHEN C=>DISPLAY<=DIG3;
        IF (PARO='0') THEN
            EDO_FUT<=D;
        ELSE
            EDO_FUT<=C;
        END IF;

WHEN D=>DISPLAY<=DIG4;
        IF (PARO='0') THEN
            EDO_FUT<=E;
        ELSE
            EDO_FUT<=D;
        END IF;

WHEN E=>DISPLAY<=DIG5;
        IF (PARO='0') THEN
            EDO_FUT<=F;
        ELSE
            EDO_FUT<=E;
        END IF;

WHEN F=>DISPLAY<=DIG6;
        IF (PARO='0') THEN
            EDO_FUT<=A;
        ELSE
            EDO_FUT<=F;
        END IF;

WHEN APAGADO=>DISPLAY <= "1111111";
                IF PARO = '0' THEN
                    EDO_FUT <= A;
                ELSE
                    EDO_FUT <= APAGADO;
                END IF;
END CASE;
END PROCESS;
PROCESS(CLR,DIV_CLK) IS
    BEGIN
    IF(CLR='0')THEN
        EDO_PRE<=APAGADO;
    ELSIF RISING_EDGE(DIV_CLK)THEN
        EDO_PRE<= EDO_FUT;
    END IF;
END PROCESS;

END ARCHITECTURE A_DADO;
